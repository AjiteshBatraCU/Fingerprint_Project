// prj_processor.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module prj_processor (
		input  wire [1:0] buttons_external_connection_export,  //  buttons_external_connection.export
		input  wire       clk_clk,                             //                          clk.clk
		input  wire       fp1_rxd,                             //                          fp1.rxd
		output wire       fp1_txd,                             //                             .txd
		input  wire       fp2_rxd,                             //                          fp2.rxd
		output wire       fp2_txd,                             //                             .txd
		output wire [7:0] hex_0_external_connection_export,    //    hex_0_external_connection.export
		output wire [7:0] hex_1_external_connection_export,    //    hex_1_external_connection.export
		output wire [7:0] hex_2_external_connection_export,    //    hex_2_external_connection.export
		output wire [7:0] hex_3_external_connection_export,    //    hex_3_external_connection.export
		output wire [7:0] hex_4_external_connection_export,    //    hex_4_external_connection.export
		output wire [7:0] hex_5_external_connection_export,    //    hex_5_external_connection.export
		output wire [9:0] leds_external_connection_export,     //     leds_external_connection.export
		output wire [7:0] pwm_control_export,                  //                  pwm_control.export
		input  wire       reset_reset_n,                       //                        reset.reset_n
		input  wire [8:0] switches_external_connection_export  // switches_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [18:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [18:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_pwm_control_s1_chipselect;               // mm_interconnect_0:PWM_control_s1_chipselect -> PWM_control:chipselect
	wire  [31:0] mm_interconnect_0_pwm_control_s1_readdata;                 // PWM_control:readdata -> mm_interconnect_0:PWM_control_s1_readdata
	wire   [1:0] mm_interconnect_0_pwm_control_s1_address;                  // mm_interconnect_0:PWM_control_s1_address -> PWM_control:address
	wire         mm_interconnect_0_pwm_control_s1_write;                    // mm_interconnect_0:PWM_control_s1_write -> PWM_control:write_n
	wire  [31:0] mm_interconnect_0_pwm_control_s1_writedata;                // mm_interconnect_0:PWM_control_s1_writedata -> PWM_control:writedata
	wire         mm_interconnect_0_fp1_control_s1_chipselect;               // mm_interconnect_0:fp1_control_s1_chipselect -> fp1_control:chipselect
	wire  [15:0] mm_interconnect_0_fp1_control_s1_readdata;                 // fp1_control:readdata -> mm_interconnect_0:fp1_control_s1_readdata
	wire   [2:0] mm_interconnect_0_fp1_control_s1_address;                  // mm_interconnect_0:fp1_control_s1_address -> fp1_control:address
	wire         mm_interconnect_0_fp1_control_s1_read;                     // mm_interconnect_0:fp1_control_s1_read -> fp1_control:read_n
	wire         mm_interconnect_0_fp1_control_s1_begintransfer;            // mm_interconnect_0:fp1_control_s1_begintransfer -> fp1_control:begintransfer
	wire         mm_interconnect_0_fp1_control_s1_write;                    // mm_interconnect_0:fp1_control_s1_write -> fp1_control:write_n
	wire  [15:0] mm_interconnect_0_fp1_control_s1_writedata;                // mm_interconnect_0:fp1_control_s1_writedata -> fp1_control:writedata
	wire         mm_interconnect_0_fp2_control_s1_chipselect;               // mm_interconnect_0:fp2_control_s1_chipselect -> fp2_control:chipselect
	wire  [15:0] mm_interconnect_0_fp2_control_s1_readdata;                 // fp2_control:readdata -> mm_interconnect_0:fp2_control_s1_readdata
	wire   [2:0] mm_interconnect_0_fp2_control_s1_address;                  // mm_interconnect_0:fp2_control_s1_address -> fp2_control:address
	wire         mm_interconnect_0_fp2_control_s1_read;                     // mm_interconnect_0:fp2_control_s1_read -> fp2_control:read_n
	wire         mm_interconnect_0_fp2_control_s1_begintransfer;            // mm_interconnect_0:fp2_control_s1_begintransfer -> fp2_control:begintransfer
	wire         mm_interconnect_0_fp2_control_s1_write;                    // mm_interconnect_0:fp2_control_s1_write -> fp2_control:write_n
	wire  [15:0] mm_interconnect_0_fp2_control_s1_writedata;                // mm_interconnect_0:fp2_control_s1_writedata -> fp2_control:writedata
	wire         mm_interconnect_0_prog_mem_s1_chipselect;                  // mm_interconnect_0:prog_mem_s1_chipselect -> prog_mem:chipselect
	wire  [31:0] mm_interconnect_0_prog_mem_s1_readdata;                    // prog_mem:readdata -> mm_interconnect_0:prog_mem_s1_readdata
	wire  [14:0] mm_interconnect_0_prog_mem_s1_address;                     // mm_interconnect_0:prog_mem_s1_address -> prog_mem:address
	wire   [3:0] mm_interconnect_0_prog_mem_s1_byteenable;                  // mm_interconnect_0:prog_mem_s1_byteenable -> prog_mem:byteenable
	wire         mm_interconnect_0_prog_mem_s1_write;                       // mm_interconnect_0:prog_mem_s1_write -> prog_mem:write
	wire  [31:0] mm_interconnect_0_prog_mem_s1_writedata;                   // mm_interconnect_0:prog_mem_s1_writedata -> prog_mem:writedata
	wire         mm_interconnect_0_prog_mem_s1_clken;                       // mm_interconnect_0:prog_mem_s1_clken -> prog_mem:clken
	wire         mm_interconnect_0_sys_timer_s1_chipselect;                 // mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_timer_s1_readdata;                   // sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_timer_s1_address;                    // mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_0_sys_timer_s1_write;                      // mm_interconnect_0:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_timer_s1_writedata;                  // mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                     // mm_interconnect_0:HEX_5_s1_chipselect -> HEX_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                       // HEX_5:readdata -> mm_interconnect_0:HEX_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                        // mm_interconnect_0:HEX_5_s1_address -> HEX_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                          // mm_interconnect_0:HEX_5_s1_write -> HEX_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                      // mm_interconnect_0:HEX_5_s1_writedata -> HEX_5:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                     // mm_interconnect_0:HEX_4_s1_chipselect -> HEX_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                       // HEX_4:readdata -> mm_interconnect_0:HEX_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                        // mm_interconnect_0:HEX_4_s1_address -> HEX_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                          // mm_interconnect_0:HEX_4_s1_write -> HEX_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                      // mm_interconnect_0:HEX_4_s1_writedata -> HEX_4:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                     // mm_interconnect_0:HEX_0_s1_chipselect -> HEX_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                       // HEX_0:readdata -> mm_interconnect_0:HEX_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                        // mm_interconnect_0:HEX_0_s1_address -> HEX_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                          // mm_interconnect_0:HEX_0_s1_write -> HEX_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                      // mm_interconnect_0:HEX_0_s1_writedata -> HEX_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                     // mm_interconnect_0:HEX_1_s1_chipselect -> HEX_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                       // HEX_1:readdata -> mm_interconnect_0:HEX_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                        // mm_interconnect_0:HEX_1_s1_address -> HEX_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                          // mm_interconnect_0:HEX_1_s1_write -> HEX_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                      // mm_interconnect_0:HEX_1_s1_writedata -> HEX_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                     // mm_interconnect_0:HEX_2_s1_chipselect -> HEX_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                       // HEX_2:readdata -> mm_interconnect_0:HEX_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                        // mm_interconnect_0:HEX_2_s1_address -> HEX_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                          // mm_interconnect_0:HEX_2_s1_write -> HEX_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                      // mm_interconnect_0:HEX_2_s1_writedata -> HEX_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                     // mm_interconnect_0:HEX_3_s1_chipselect -> HEX_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                       // HEX_3:readdata -> mm_interconnect_0:HEX_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                        // mm_interconnect_0:HEX_3_s1_address -> HEX_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                          // mm_interconnect_0:HEX_3_s1_write -> HEX_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                      // mm_interconnect_0:HEX_3_s1_writedata -> HEX_3:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                      // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                        // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                         // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                           // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                       // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                     // Buttons:readdata -> mm_interconnect_0:Buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                      // mm_interconnect_0:Buttons_s1_address -> Buttons:address
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                    // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                     // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire         irq_mapper_receiver0_irq;                                  // fp1_control:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // fp2_control:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // sys_timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [Buttons:reset_n, HEX_0:reset_n, HEX_1:reset_n, HEX_2:reset_n, HEX_3:reset_n, HEX_4:reset_n, HEX_5:reset_n, LEDs:reset_n, PWM_control:reset_n, Switches:reset_n, cpu:reset_n, fp1_control:reset_n, fp2_control:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, prog_mem:reset, rst_translator:in_reset, sys_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, prog_mem:reset_req, rst_translator:reset_req_in]

	prj_processor_Buttons buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_external_connection_export)     // external_connection.export
	);

	prj_processor_HEX_0 hex_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex_0_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 hex_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex_1_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 hex_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex_2_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 hex_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex_3_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 hex_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex_4_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 hex_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex_5_external_connection_export)       // external_connection.export
	);

	prj_processor_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	prj_processor_HEX_0 pwm_control (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pwm_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm_control_s1_readdata),   //                    .readdata
		.out_port   (pwm_control_export)                           // external_connection.export
	);

	prj_processor_Switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	prj_processor_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	prj_processor_fp1_control fp1_control (
		.clk           (clk_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address       (mm_interconnect_0_fp1_control_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_fp1_control_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_fp1_control_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_fp1_control_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_fp1_control_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_fp1_control_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_fp1_control_s1_readdata),      //                    .readdata
		.rxd           (fp1_rxd),                                        // external_connection.export
		.txd           (fp1_txd),                                        //                    .export
		.irq           (irq_mapper_receiver0_irq)                        //                 irq.irq
	);

	prj_processor_fp1_control fp2_control (
		.clk           (clk_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address       (mm_interconnect_0_fp2_control_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_fp2_control_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_fp2_control_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_fp2_control_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_fp2_control_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_fp2_control_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_fp2_control_s1_readdata),      //                    .readdata
		.rxd           (fp2_rxd),                                        // external_connection.export
		.txd           (fp2_txd),                                        //                    .export
		.irq           (irq_mapper_receiver1_irq)                        //                 irq.irq
	);

	prj_processor_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	prj_processor_prog_mem prog_mem (
		.clk        (clk_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_prog_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_prog_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_prog_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_prog_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_prog_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_prog_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_prog_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	prj_processor_sys_timer sys_timer (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                   //   irq.irq
	);

	prj_processor_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	prj_processor_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                         clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_readdatavalid           (cpu_data_master_readdatavalid),                             //                                .readdatavalid
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                .readdatavalid
		.Buttons_s1_address                      (mm_interconnect_0_buttons_s1_address),                      //                      Buttons_s1.address
		.Buttons_s1_readdata                     (mm_interconnect_0_buttons_s1_readdata),                     //                                .readdata
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.fp1_control_s1_address                  (mm_interconnect_0_fp1_control_s1_address),                  //                  fp1_control_s1.address
		.fp1_control_s1_write                    (mm_interconnect_0_fp1_control_s1_write),                    //                                .write
		.fp1_control_s1_read                     (mm_interconnect_0_fp1_control_s1_read),                     //                                .read
		.fp1_control_s1_readdata                 (mm_interconnect_0_fp1_control_s1_readdata),                 //                                .readdata
		.fp1_control_s1_writedata                (mm_interconnect_0_fp1_control_s1_writedata),                //                                .writedata
		.fp1_control_s1_begintransfer            (mm_interconnect_0_fp1_control_s1_begintransfer),            //                                .begintransfer
		.fp1_control_s1_chipselect               (mm_interconnect_0_fp1_control_s1_chipselect),               //                                .chipselect
		.fp2_control_s1_address                  (mm_interconnect_0_fp2_control_s1_address),                  //                  fp2_control_s1.address
		.fp2_control_s1_write                    (mm_interconnect_0_fp2_control_s1_write),                    //                                .write
		.fp2_control_s1_read                     (mm_interconnect_0_fp2_control_s1_read),                     //                                .read
		.fp2_control_s1_readdata                 (mm_interconnect_0_fp2_control_s1_readdata),                 //                                .readdata
		.fp2_control_s1_writedata                (mm_interconnect_0_fp2_control_s1_writedata),                //                                .writedata
		.fp2_control_s1_begintransfer            (mm_interconnect_0_fp2_control_s1_begintransfer),            //                                .begintransfer
		.fp2_control_s1_chipselect               (mm_interconnect_0_fp2_control_s1_chipselect),               //                                .chipselect
		.HEX_0_s1_address                        (mm_interconnect_0_hex_0_s1_address),                        //                        HEX_0_s1.address
		.HEX_0_s1_write                          (mm_interconnect_0_hex_0_s1_write),                          //                                .write
		.HEX_0_s1_readdata                       (mm_interconnect_0_hex_0_s1_readdata),                       //                                .readdata
		.HEX_0_s1_writedata                      (mm_interconnect_0_hex_0_s1_writedata),                      //                                .writedata
		.HEX_0_s1_chipselect                     (mm_interconnect_0_hex_0_s1_chipselect),                     //                                .chipselect
		.HEX_1_s1_address                        (mm_interconnect_0_hex_1_s1_address),                        //                        HEX_1_s1.address
		.HEX_1_s1_write                          (mm_interconnect_0_hex_1_s1_write),                          //                                .write
		.HEX_1_s1_readdata                       (mm_interconnect_0_hex_1_s1_readdata),                       //                                .readdata
		.HEX_1_s1_writedata                      (mm_interconnect_0_hex_1_s1_writedata),                      //                                .writedata
		.HEX_1_s1_chipselect                     (mm_interconnect_0_hex_1_s1_chipselect),                     //                                .chipselect
		.HEX_2_s1_address                        (mm_interconnect_0_hex_2_s1_address),                        //                        HEX_2_s1.address
		.HEX_2_s1_write                          (mm_interconnect_0_hex_2_s1_write),                          //                                .write
		.HEX_2_s1_readdata                       (mm_interconnect_0_hex_2_s1_readdata),                       //                                .readdata
		.HEX_2_s1_writedata                      (mm_interconnect_0_hex_2_s1_writedata),                      //                                .writedata
		.HEX_2_s1_chipselect                     (mm_interconnect_0_hex_2_s1_chipselect),                     //                                .chipselect
		.HEX_3_s1_address                        (mm_interconnect_0_hex_3_s1_address),                        //                        HEX_3_s1.address
		.HEX_3_s1_write                          (mm_interconnect_0_hex_3_s1_write),                          //                                .write
		.HEX_3_s1_readdata                       (mm_interconnect_0_hex_3_s1_readdata),                       //                                .readdata
		.HEX_3_s1_writedata                      (mm_interconnect_0_hex_3_s1_writedata),                      //                                .writedata
		.HEX_3_s1_chipselect                     (mm_interconnect_0_hex_3_s1_chipselect),                     //                                .chipselect
		.HEX_4_s1_address                        (mm_interconnect_0_hex_4_s1_address),                        //                        HEX_4_s1.address
		.HEX_4_s1_write                          (mm_interconnect_0_hex_4_s1_write),                          //                                .write
		.HEX_4_s1_readdata                       (mm_interconnect_0_hex_4_s1_readdata),                       //                                .readdata
		.HEX_4_s1_writedata                      (mm_interconnect_0_hex_4_s1_writedata),                      //                                .writedata
		.HEX_4_s1_chipselect                     (mm_interconnect_0_hex_4_s1_chipselect),                     //                                .chipselect
		.HEX_5_s1_address                        (mm_interconnect_0_hex_5_s1_address),                        //                        HEX_5_s1.address
		.HEX_5_s1_write                          (mm_interconnect_0_hex_5_s1_write),                          //                                .write
		.HEX_5_s1_readdata                       (mm_interconnect_0_hex_5_s1_readdata),                       //                                .readdata
		.HEX_5_s1_writedata                      (mm_interconnect_0_hex_5_s1_writedata),                      //                                .writedata
		.HEX_5_s1_chipselect                     (mm_interconnect_0_hex_5_s1_chipselect),                     //                                .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.LEDs_s1_address                         (mm_interconnect_0_leds_s1_address),                         //                         LEDs_s1.address
		.LEDs_s1_write                           (mm_interconnect_0_leds_s1_write),                           //                                .write
		.LEDs_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                        //                                .readdata
		.LEDs_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                       //                                .writedata
		.LEDs_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                      //                                .chipselect
		.prog_mem_s1_address                     (mm_interconnect_0_prog_mem_s1_address),                     //                     prog_mem_s1.address
		.prog_mem_s1_write                       (mm_interconnect_0_prog_mem_s1_write),                       //                                .write
		.prog_mem_s1_readdata                    (mm_interconnect_0_prog_mem_s1_readdata),                    //                                .readdata
		.prog_mem_s1_writedata                   (mm_interconnect_0_prog_mem_s1_writedata),                   //                                .writedata
		.prog_mem_s1_byteenable                  (mm_interconnect_0_prog_mem_s1_byteenable),                  //                                .byteenable
		.prog_mem_s1_chipselect                  (mm_interconnect_0_prog_mem_s1_chipselect),                  //                                .chipselect
		.prog_mem_s1_clken                       (mm_interconnect_0_prog_mem_s1_clken),                       //                                .clken
		.PWM_control_s1_address                  (mm_interconnect_0_pwm_control_s1_address),                  //                  PWM_control_s1.address
		.PWM_control_s1_write                    (mm_interconnect_0_pwm_control_s1_write),                    //                                .write
		.PWM_control_s1_readdata                 (mm_interconnect_0_pwm_control_s1_readdata),                 //                                .readdata
		.PWM_control_s1_writedata                (mm_interconnect_0_pwm_control_s1_writedata),                //                                .writedata
		.PWM_control_s1_chipselect               (mm_interconnect_0_pwm_control_s1_chipselect),               //                                .chipselect
		.Switches_s1_address                     (mm_interconnect_0_switches_s1_address),                     //                     Switches_s1.address
		.Switches_s1_readdata                    (mm_interconnect_0_switches_s1_readdata),                    //                                .readdata
		.sys_timer_s1_address                    (mm_interconnect_0_sys_timer_s1_address),                    //                    sys_timer_s1.address
		.sys_timer_s1_write                      (mm_interconnect_0_sys_timer_s1_write),                      //                                .write
		.sys_timer_s1_readdata                   (mm_interconnect_0_sys_timer_s1_readdata),                   //                                .readdata
		.sys_timer_s1_writedata                  (mm_interconnect_0_sys_timer_s1_writedata),                  //                                .writedata
		.sys_timer_s1_chipselect                 (mm_interconnect_0_sys_timer_s1_chipselect),                 //                                .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //             sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata)             //                                .readdata
	);

	prj_processor_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
